ENTITY A IS

END ENTITY A;