PACKAGE n IS -- This is a comment
END PACKAGE n;